module TimeDisplayMode(
    input sw,
    input TSmode_state,
    input SSmode_state,
    output TDmode_state
);
// 각각의 모드에서 어떤 state인가에 따라서 TDmode 내 state 이동을 결정한다


endmodule

